module andgate_df(a,b,y);
input a,b;
output y;
  assign y=a&b;  //and(y,a,b)
endmodule
